
package mypackage is

	type ImageMatrix is array(natural range <>, natural range <>) of std_logic_vector(23 downto 0);

	type KernalMatrix is array(natural range <>, natural range <>) of std_logic_vector(7 downto 0);

end package mypackage;

